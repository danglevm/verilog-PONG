module UART_RX (

);